module {name}_core;
endmodule
