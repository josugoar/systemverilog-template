package {name}_pkg;
endpackage
